localparam ccd_mode_idle        = 2'b00;
localparam ccd_mode_clean       = 2'b01;
localparam ccd_mode_readout_1x1 = 2'b10;
localparam ccd_mode_readout_2x2 = 2'b11;
